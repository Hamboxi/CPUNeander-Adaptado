library verilog;
use verilog.vl_types.all;
entity PEx03SomadorSubtradorAcumulador_vlg_vec_tst is
end PEx03SomadorSubtradorAcumulador_vlg_vec_tst;
