library verilog;
use verilog.vl_types.all;
entity MEM_vlg_vec_tst is
end MEM_vlg_vec_tst;
